-------------------------------------------------------------------------------
--
-- CDC 6600 model
--
-- Copyright (C) 2010 by Paul Koning
--
-- Derived from the original 6600 module design
-- by Seymour Cray and his team at Control Data,
-- as documented in CDC 6600 "Chassis Tabs" manuals,
-- which are in the public domain.  Scans supplied
-- from the Computer History Museum collection
-- by Dave Redell and Al Kossow.
--
-- TP module
--
-------------------------------------------------------------------------------

use work.sigs.all;

entity tp is
    port (
      p1 : in  logicsig;
      p13 : in  logicsig;
      p14 : in  logicsig;
      p15 : in  logicsig;
      p27 : in  logicsig;
      p28 : in  logicsig;
      tp1 : out logicsig;
      tp2 : out logicsig;
      tp3 : out logicsig;
      tp4 : out logicsig;
      tp5 : out logicsig;
      tp6 : out logicsig;
      p2 : out logicsig;
      p3 : out logicsig;
      p4 : out logicsig;
      p5 : out logicsig;
      p6 : out logicsig;
      p7 : out logicsig;
      p8 : out logicsig;
      p9 : out logicsig;
      p10 : out logicsig;
      p11 : out logicsig;
      p12 : out logicsig;
      p16 : out logicsig;
      p17 : out logicsig;
      p18 : out logicsig;
      p19 : out logicsig;
      p20 : out logicsig;
      p21 : out logicsig;
      p22 : out logicsig;
      p23 : out logicsig;
      p24 : out logicsig;
      p25 : out logicsig;
      p26 : out logicsig);

end tp;
architecture gates of tp is
  component g2
    port (
      a : in  logicsig;
      b : in  logicsig;
      y : out logicsig;
      y2 : out logicsig);

  end component;

  component inv2
    port (
      a : in  logicsig;
      y : out logicsig;
      y2 : out logicsig);

  end component;

  signal t1 : logicsig;
  signal t2 : logicsig;
  signal t3 : logicsig;
  signal t4 : logicsig;

begin -- gates
  u1 : inv2 port map (
    a => p1,
    y => tp1,
    y2 => t1);

  p3 <= t1;
  p5 <= t1;
  p7 <= t1;
  p9 <= t1;
  p11 <= t1;

  u2 : inv2 port map (
    a => p14,
    y => tp2,
    y2 => t2);

  p2 <= t2;
  p4 <= t2;
  p6 <= t2;
  p8 <= t2;
  p10 <= t2;
  p12 <= t2;
  tp3 <= t2;

  u3 : g2 port map (
    a => p13,
    b => p15,
    y => tp4,
    y2 => t3);

  p17 <= t3;
  p19 <= t3;
  p21 <= t3;
  p23 <= t3;
  p25 <= t3;

  u4 : g2 port map (
    a => p27,
    b => p28,
    y => tp5,
    y2 => t4);

  p16 <= t4;
  p18 <= t4;
  p20 <= t4;
  p22 <= t4;
  p24 <= t4;
  p26 <= t4;
  tp6 <= t4;


end gates;

