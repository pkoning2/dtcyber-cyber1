-------------------------------------------------------------------------------
--
-- CDC 6600 model
--
-- Copyright (C) 2009 by Paul Koning
--
-- Derived from the original 6600 module design
-- by Seymour Cray and his team at Control Data,
-- as documented in CDC 6600 "Chassis Tabs" manuals,
-- which are in the public domain.  Scans supplied
-- from the Computer History Museum collection
-- by Dave Redell and Al Kossow.
--
-- HB module
--
-------------------------------------------------------------------------------

use work.sigs.all;

entity hb is
    port (
      p13 : in  logicsig;
      p14 : in  logicsig;
      p15 : in  logicsig;
      p16 : in  logicsig;
      tp1 : out logicsig;
      tp2 : out logicsig;
      tp5 : out logicsig;
      tp6 : out logicsig;
      p1 : out logicsig;
      p2 : out logicsig;
      p3 : out logicsig;
      p4 : out logicsig;
      p5 : out logicsig;
      p6 : out logicsig;
      p7 : out logicsig;
      p8 : out logicsig;
      p9 : out logicsig;
      p10 : out logicsig;
      p11 : out logicsig;
      p12 : out logicsig;
      p17 : out logicsig;
      p18 : out logicsig;
      p19 : out logicsig;
      p20 : out logicsig;
      p21 : out logicsig;
      p22 : out logicsig;
      p23 : out logicsig;
      p24 : out logicsig;
      p25 : out logicsig;
      p26 : out logicsig;
      p27 : out logicsig;
      p28 : out logicsig);

end hb;
architecture gates of hb is
  component g2
    port (
      a : in  logicsig;
      b : in  logicsig;
      y : out logicsig;
      y2 : out logicsig);

  end component;

  component inv2
    port (
      a : in  logicsig;
      y : out logicsig;
      y2 : out logicsig);

  end component;

  signal t1 : logicsig;
  signal t2 : logicsig;
  signal t3 : logicsig;
  signal t4 : logicsig;
  signal t5 : logicsig;
  signal t6 : logicsig;
  signal t7 : logicsig;
  signal t8 : logicsig;

begin -- gates
  u1 : g2 port map (
    a => p13,
    b => p14,
    y2 => t1);

  p12 <= t1;
  tp1 <= t1;

  u2 : g2 port map (
    a => p14,
    b => p16,
    y2 => t2);

  p11 <= t2;
  tp2 <= t2;

  u3 : g2 port map (
    a => p13,
    b => p15,
    y2 => t3);

  p18 <= t3;
  tp5 <= t3;

  u4 : g2 port map (
    a => p16,
    b => p15,
    y2 => t4);

  p17 <= t4;
  tp6 <= t4;

  u5 : inv2 port map (
    a => t1,
    y2 => t5);

  p2 <= t5;
  p4 <= t5;
  p6 <= t5;
  p8 <= t5;
  p10 <= t5;

  u6 : inv2 port map (
    a => t2,
    y2 => t6);

  p1 <= t6;
  p3 <= t6;
  p5 <= t6;
  p7 <= t6;
  p9 <= t6;

  u7 : inv2 port map (
    a => t3,
    y2 => t7);

  p20 <= t7;
  p22 <= t7;
  p24 <= t7;
  p26 <= t7;
  p28 <= t7;

  u8 : inv2 port map (
    a => t4,
    y2 => t8);

  p19 <= t8;
  p21 <= t8;
  p23 <= t8;
  p25 <= t8;
  p27 <= t8;


end gates;

