-------------------------------------------------------------------------------
--
-- CDC 6600 model
--
-- Copyright (C) 2009 by Paul Koning
--
-- Derived from the original 6600 module design
-- by Seymour Cray and his team at Control Data,
-- as documented in CDC 6600 "Chassis Tabs" manuals,
-- which are in the public domain.  Scans supplied
-- from the Computer History Museum collection
-- by Dave Redell and Al Kossow.
--
-- AJ module
--
-------------------------------------------------------------------------------

use work.sigs.all;

entity aj is
    port (
      p1 : in  logicsig;
      p3 : in  logicsig;
      p7 : in  logicsig;
      p8 : in  logicsig;
      p9 : in  logicsig;
      p10 : in  logicsig;
      p11 : in  logicsig;
      p18 : in  logicsig;
      p20 : in  logicsig;
      p22 : in  logicsig;
      p24 : in  logicsig;
      p26 : in  logicsig;
      p28 : in  logicsig;
      tp1 : out logicsig;
      tp2 : out logicsig;
      tp5 : out logicsig;
      tp6 : out logicsig;
      p4 : out logicsig;
      p5 : out logicsig;
      p6 : out logicsig;
      p13 : out logicsig;
      p14 : out logicsig;
      p15 : out logicsig;
      p17 : out logicsig;
      p19 : out logicsig;
      p21 : out logicsig;
      p23 : out logicsig;
      p27 : out logicsig);

end aj;
architecture gates of aj is
  component g2
    port (
      a : in  logicsig;
      b : in  logicsig;
      y : out logicsig;
      y2 : out logicsig);

  end component;

  component inv
    port (
      a : in  logicsig;
      y : out logicsig);

  end component;

  component inv2
    port (
      a : in  logicsig;
      y : out logicsig;
      y2 : out logicsig);

  end component;

  component latch22
    port (
      clk : in  logicsig;
      clk2 : in  logicsig;
      d : in  logicsig;
      d2 : in  logicsig;
      q : out logicsig;
      qb : out logicsig);

  end component;

  component rs2flop
    port (
      r : in  logicsig;
      s : in  logicsig;
      s2 : in  logicsig;
      q : out logicsig;
      qb : out logicsig);

  end component;

  signal a : logicsig;
  signal b : logicsig;
  signal t2 : logicsig;
  signal t4 : logicsig;
  signal t7 : logicsig;
  signal t8 : logicsig;
  signal t11 : logicsig;
  signal t12 : logicsig;

begin -- gates
  u2 : g2 port map (
    a => p1,
    b => p3,
    y => t2);

  u3 : latch22 port map (
    clk  => p7,
    clk2 => p22,
    d    => a,
    d2   => t2,
    q    => t4);

  p4 <= t4;
  tp1 <= t4;

  u5 : g2 port map (
    a => t4,
    b => p10,
    y => p6);


  u7 : g2 port map (
    a => p28,
    b => p26,
    y => t7);


  u8 : latch22 port map (
    clk  => p7,
    clk2 => p22,
    d    => b,
    d2   => t7,
    q    => t8,
    qb   => p23);

  p14 <= t8;
  p21 <= t8;
  tp6 <= t8;

  u9 : inv port map (
    a => t8,
    y => p5);

  
  u10 : g2 port map (
    a => p24,
    b => t8,
    y => p27);


  u11 : rs2flop port map (
    r => t11,
    s => p11,
    s2 => p9,
    q => a);

  tp2 <= a;


  u13 : inv2 port map (
    a => p8,
    y => t11,
    y2 => t12);

  p13 <= t12;
  p15 <= t12;
  p17 <= t12;
  p19 <= t12;

  u14 : rs2flop port map (
    r => t11,
    s => p20,
    s2 => p18,
    q => b);

  tp5 <= b;


end gates;

